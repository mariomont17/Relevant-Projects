package params_pkg;
  parameter TERMINALES = 10;
  parameter PROFUNDIDAD = 31;
endpackage
