package params_pkg;
  parameter PROFUNDIDAD = 30;
endpackage